library verilog;
use verilog.vl_types.all;
entity TL_vlg_vec_tst is
end TL_vlg_vec_tst;
