library verilog;
use verilog.vl_types.all;
entity prueba_vlg_vec_tst is
end prueba_vlg_vec_tst;
